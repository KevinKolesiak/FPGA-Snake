// Snake Game interface
// Kevin Kolesiak

//instantiate balls to be appended to 

//head ball


//module game_interface ( input Reset, frame_clk, input [7:0] keycode, 
//								output [9:0]  BallX, BallY, BallS, FoodX, FoodY, FoodS);
//
//



//ball Head(.Reset(Reset_h), .frame_clk(VGA_VS), .keycode(keycode),
//               .BallX(ballxsig), .BallY(ballysig), .BallS(ballsizesig)
//);


//all other balls



//instantiate food in random positions


//endmodule
